module alu #(parameter OPSIZE = 4, parameter DSIZE = 16)(
  output [DSIZE-1:0] F
);

endmodule